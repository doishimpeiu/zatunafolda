module w1 (
  output [3:0] w0_raddr,
  input signed [7:0] w0_rdata,
  output [3:0] w1_raddr,
  input signed [7:0] w1_rdata,
  output [3:0] w2_raddr,
  input signed [7:0] w2_rdata,
  output [3:0] w3_raddr,
  input signed [7:0] w3_rdata,
  output [3:0] w4_raddr,
  input signed [7:0] w4_rdata,
  output [3:0] w5_raddr,
  input signed [7:0] w5_rdata,
  output [3:0] w6_raddr,
  input signed [7:0] w6_rdata,
  output [3:0] w7_raddr,
  input signed [7:0] w7_rdata,
  output [3:0] w8_raddr,
  input signed [7:0] w8_rdata,
  output [3:0] w9_raddr,
  input signed [7:0] w9_rdata,
  output [3:0] w10_raddr,
  input signed [7:0] w10_rdata,
  output [3:0] w11_raddr,
  input signed [7:0] w11_rdata,
  output [3:0] w12_raddr,
  input signed [7:0] w12_rdata,
  output [3:0] w13_raddr,
  input signed [7:0] w13_rdata,
  output [3:0] w14_raddr,
  input signed [7:0] w14_rdata,
  output [3:0] w15_raddr,
  input signed [7:0] w15_rdata,
  input start,
  output finish,
  input clk, xrst
);